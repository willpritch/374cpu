module DataPath(
	input wire clock, clear,
	input wire [31:0] Mdatain,
	input wire [4:0] opcode,
	
	input RAout, R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out, 
	RYout, RZHIout, RZLOout, PCout, IRout, HIout, LOout, MDRout, PORTout,
	
	input RAin, R0in, R1in, R2in, R3in, R4in, R5in, R6in, R7in, R8in, R9in, R10in, R11in, R12in, R13in, R14in, R15in, 
	RYin, RZin, PCin, IRin, HIin, LOin, MDRin, PORTin, Read
	
	);

wire [31:0] BusMuxOut, BusMuxInRA, BusMuxInR0, BusMuxInR1, BusMuxInR2, BusMuxInR3, BusMuxInR4, BusMuxInR5, BusMuxInR6, BusMuxInR7, BusMuxInR8, 
	BusMuxInR9, BusMuxInR10, BusMuxInR11,BusMuxInR12, BusMuxInR13, BusMuxInR14, BusMuxInR15, RYdataout, BusMuxInHI, BusMuxInLO, BusMuxInRZHI, BusMuxInRZLO, 
	BusMuxInPC, BusMuxInMDR, BusMuxInPort, BusMuxInIR, RegisterAImmediate;
	
wire [63:0] Zin;

REG RA(clear, clock, RAin, RegisterAImmediate, BusMuxInRA);

REG R0(clear, clock, R0in, BusMuxOut, BusMuxInR0);
REG R1(clear, clock, R1in, BusMuxOut, BusMuxInR1);
REG R2(clear, clock, R2in, BusMuxOut, BusMuxInR2);
REG R3(clear, clock, R3in, BusMuxOut, BusMuxInR3);
REG R4(clear, clock, R4in, BusMuxOut, BusMuxInR4);
REG R5(clear, clock, R5in, BusMuxOut, BusMuxInR5);
REG R6(clear, clock, R6in, BusMuxOut, BusMuxInR6);
REG R7(clear, clock, R7in, BusMuxOut, BusMuxInR7);
REG R8(clear, clock, R8in, BusMuxOut, BusMuxInR8);	
REG R9(clear, clock, R9in, BusMuxOut, BusMuxInR9);
REG R10(clear, clock, R10in, BusMuxOut, BusMuxInR10);
REG R11(clear, clock, R11in, BusMuxOut, BusMuxInR11);
REG R12(clear, clock, R12in, BusMuxOut, BusMuxInR12);
REG R13(clear, clock, R13in, BusMuxOut, BusMuxInR13);
REG R14(clear, clock, R14in, BusMuxOut, BusMuxInR14);
REG R15(clear, clock, R15in, BusMuxOut, BusMuxInR15);
REG RY(clear, clock, RYin, BusMuxOut, RYdataout);
REG RZHI(clear, clock, RZin, Zin[63:32], BusMuxInRZHI); 
REG RZLO(clear, clock, RZin, Zin[31:0], BusMuxInRZLO); 
REG PC(clear, clock, PCin, BusMuxOut, BusMuxInPC);
REG IR(clear, clock, IRin, BusMuxOut, BusMuxInIR);
REG HI(clear, clock, HIin, BusMuxOut, BusMuxInHI);
REG LO(clear, clock, LOin, BusMuxOut, BusMuxInLO);

Bus bus(BusMuxInRA, BusMuxInR0, BusMuxInR1, BusMuxInR2, BusMuxInR3, BusMuxInR4, BusMuxInR5, BusMuxInR6, BusMuxInR7, BusMuxInR8, 
	BusMuxInR9, BusMuxInR10, BusMuxInR11,BusMuxInR12, BusMuxInR13, BusMuxInR14, BusMuxInR15, BusMuxInHI, BusMuxInLO, BusMuxInRZHI, BusMuxInRZLO, 
	BusMuxInPC, BusMuxInMDR, BusMuxInPort, RAout, R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, 
	R13out, R14out, R15out, RYout, RZHIout, RZLOout, PCout, IRout, HIout, LOout, MDRout, PORTout, BusMuxOut);

MDR MDR(clear, clock, MDRin, Read, Mdatain, BusMuxOut, BusMuxInMDR);

ALU ALU(opcode, RYdataout, BusMuxOut, Zin);

endmodule
